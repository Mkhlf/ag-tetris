`include "src/GLOBAL.sv"

module game_top(
    input  wire logic CLK100MHZ,
    input  wire logic CPU_RESETN, // Active Low
    input  wire logic PS2_CLK,
    input  wire logic PS2_DATA,
    input  wire logic btn_l,
    input  wire logic btn_r,
    input  wire logic btn_u,
    input  wire logic btn_d,
    input  wire logic btn_c,
    output logic [3:0] VGA_R,
    output logic [3:0] VGA_G,
    output logic [3:0] VGA_B,
    output logic VGA_HS,
    output logic VGA_VS
    );

    logic rst;
    assign rst = ~CPU_RESETN;

    // Clock Generation
    logic pix_clk; // 83.46 MHz (approx)
    logic locked;
    
    // Instantiate Clock Wizard
    clk_wiz_0 clk_gen (
        .clk_in1(CLK100MHZ),
        .clk_out1(pix_clk),
        .reset(rst),
        .locked(locked)
    );

    // Game Clock Generation (25 MHz)
    // Divide 100MHz by 4
    logic [1:0] clk_div;
    logic game_clk;
    
    always_ff @(posedge CLK100MHZ) begin
        if (rst) clk_div <= 0;
        else clk_div <= clk_div + 1;
    end
    assign game_clk = clk_div[1]; // 25 MHz

    // Game Tick Generation (60Hz)
    // 25 MHz / 60 Hz ~= 416,666
    logic [18:0] tick_counter;
    logic tick_game;
    
    always_ff @(posedge game_clk) begin
        if (rst) begin
            tick_counter <= 0;
            tick_game <= 0;
        end else begin
            if (tick_counter == 416666) begin
                tick_counter <= 0;
                tick_game <= 1;
            end else begin
                tick_counter <= tick_counter + 1;
                tick_game <= 0;
            end
        end
    end

    // Keyboard Input
    logic [7:0] scan_code;
    logic make_break;
    
    ps2_keyboard kb_inst (
        .clk(game_clk),
        .rst(rst),
        .ps2_clk(PS2_CLK),
        .ps2_data(PS2_DATA),
        .current_scan_code(scan_code),
        .current_make_break(make_break)
    );
    
    // Input Synchronizers (Robust State Machines)
    logic key_left_ps2, key_right_ps2, key_down_ps2, key_rotate_ps2, key_drop_ps2;
    
    keyboard_to_1_clock #(.SCAN_CODE(`LEFT_ARROW_C))  k_left  (.clk(game_clk), .scanCode(scan_code), .makeBreak(make_break), .signal(key_left_ps2));
    keyboard_to_1_clock #(.SCAN_CODE(`RIGHT_ARROW_C)) k_right (.clk(game_clk), .scanCode(scan_code), .makeBreak(make_break), .signal(key_right_ps2));
    keyboard_to_1_clock #(.SCAN_CODE(`DOWN_ARROW_C))  k_down  (.clk(game_clk), .scanCode(scan_code), .makeBreak(make_break), .signal(key_down_ps2));
    keyboard_to_1_clock #(.SCAN_CODE(`UP_ARROW_C))    k_up    (.clk(game_clk), .scanCode(scan_code), .makeBreak(make_break), .signal(key_rotate_ps2));
    keyboard_to_1_clock #(.SCAN_CODE(`SPACE_C))       k_space (.clk(game_clk), .scanCode(scan_code), .makeBreak(make_break), .signal(key_drop_ps2));
    
    // Combine Inputs (Buttons + Keyboard)
    logic key_left, key_right, key_down, key_rotate, key_drop;
    
    // Note: Buttons are active high. We might want to debounce them too, 
    // but for now direct ORing is fine if buttons are clean enough.
    // Ideally we'd run buttons through a synchronizer too.
    
    assign key_left   = key_left_ps2   | btn_l;
    assign key_right  = key_right_ps2  | btn_r;
    assign key_down   = key_down_ps2   | btn_d;
    assign key_rotate = key_rotate_ps2 | btn_u;
    assign key_drop   = key_drop_ps2   | btn_c;

    // Game Logic
    field_t display_field;
    logic [31:0] score;
    logic game_over;
    
    game_control game_inst (
        .clk(game_clk),
        .rst(rst),
        .tick_game(tick_game),
        .key_left(key_left),
        .key_right(key_right),
        .key_down(key_down),
        .key_rotate(key_rotate),
        .key_drop(key_drop),
        .display(display_field),
        .score(score),
        .game_over(game_over)
    );

    // VGA Output (Raw)
    logic [10:0] curr_x_raw;
    logic [9:0]  curr_y_raw;
    logic active_area_raw;
    logic hsync_raw, vsync_raw;
    
    vga_out vga_inst (
        .clk(pix_clk),
        .rst(rst),
        .curr_x(curr_x_raw),
        .curr_y(curr_y_raw),
        .hsync(hsync_raw),
        .vsync(vsync_raw),
        .active_area(active_area_raw)
    );

    // Sprite ROM
    logic [3:0] sprite_addr_x;
    logic [3:0] sprite_addr_y;
    logic [11:0] sprite_pixel;
    
    block_sprite sprite_inst (
        .clk(pix_clk),
        .addr_x(sprite_addr_x),
        .addr_y(sprite_addr_y),
        .pixel_out(sprite_pixel)
    );

    // Drawing Logic (Raw)
    logic [3:0] vga_r_raw, vga_g_raw, vga_b_raw;

    draw_tetris draw_inst (
        .clk(pix_clk),
        .curr_x(curr_x_raw),
        .curr_y(curr_y_raw),
        .active_area(active_area_raw),
        .display(display_field),
        .score(score),
        .game_over(game_over),
        .sprite_addr_x(sprite_addr_x),
        .sprite_addr_y(sprite_addr_y),
        .sprite_pixel(sprite_pixel),
        .vga_r(vga_r_raw),
        .vga_g(vga_g_raw),
        .vga_b(vga_b_raw)
    );

    // Output Pipeline (Fix Ghosting)
    always_ff @(posedge pix_clk) begin
        VGA_R <= vga_r_raw;
        VGA_G <= vga_g_raw;
        VGA_B <= vga_b_raw;
        VGA_HS <= hsync_raw;
        VGA_VS <= vsync_raw;
    end

endmodule
